circuit 1 - linear

.options nobypass
.options

R1 1 0 1k
I1 1 0 dc -0.001

.print op v(1) i(R1)
.op

.end
