circuit 1

*.options dampmax=1.0
*.options dampmin=0.5

R1 1 0 1k
I1 1 0 dc -0.001

R2 1 2 5k
d3 2 0 dio1

.model dio1 d is=1.e-12

.print op v(1) v(2) i(R2)
.op

.end
