* example1
*.options parhier - not implemented in ltspice  - hspice specific
.options parhier=local

.param a='1'
.param w='5'

.subckt VOLTS n1 n2 n3 x='w'

*.param w='3'
.param b='2'
.param c='x'
v1 n1 0 'a'
v2 n2 0 'b'
v3 n3 0 'c'
.ends


.subckt VOLTS1 n1 n2 n3 x='w'

.param w='3'
.param b='2'
.param c='x'
v1 n1 0 'a'
v2 n2 0 'b'
v3 n3 0 'c'
.ends

X1 1 2 3 VOLTS
x2 4 5 6 VOLTS1

* result:
* 1 2 5 1 2 3 
* means that in subckt VOLTS1 w='3' overrides upper-level 'w'=5 _before_ execution of x='w'
* i.e. caclulation is carries in the sequence:
* compute c: c=x
* compute x: x=w
* compute w: w=3 (case of VOLTS1)
* hslice parhier-local - gives the same result
* if parhier-global - result like in VOLTS
* 1 2 5 1 2 5

.print  v(1) v(2) v(3) v(4) v(5) v(6) 
.op
.end

