* test for substitution
.options dollar_as_spice_comment
.attach ./bsim330.so

v1 n1 0 dc 1  
 
.list
.end
