circuit 1 - MAIN NOW

*.options dampmax=1.0
*.options dampmin=0.5

R1 1 0 1k
I1 1 0 dc -0.001
A3 1 0 amodel1 0.001

.model amodel1 A 

.print op v(1) i(R1)
.op

.end
