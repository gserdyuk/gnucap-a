circuit 1

V1 1 0 dc 1

R1 1 2 5k
R1 2 0 2.5k


.print op v(1) i(R1)
.op

.end
