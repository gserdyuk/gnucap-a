v2 n2 0 dc 2
 