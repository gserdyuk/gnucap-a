* test for substitution
#.options dollar_as_spice_comment
#.options

v1 n1 0 dc 1  
.include $PWD2/lib_file2.ckt
 
.list
.print op v(n*)
.op
.end
