v3 n3 0 dc 3
 