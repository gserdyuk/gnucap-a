noise - sources manipulation + - - 
v1   1  0  dc 1 ac 1
R1   1  0  100.
R2   1  2  10
R3   2  0  100


.print noise inoise
.print noise + onoise
.print noise - inoise onoise
.noise v(2) v1 dec 10 10 100

.end
