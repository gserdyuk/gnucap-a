v4 n4 0 dc 4
 