circuit 1

R1 1 0 1k
I1 1 0 dc 0.001

R2 1 2 5k
R3 2 0 2.5k

.print op v(1) i(R1)
.op

.end
