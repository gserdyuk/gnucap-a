circuit 2 - cubic

.options nobypass
*.options

A1 1 0 deva1 AR=0.001 B=0.001 V0=1
I1 1 0 dc -0.001

.model deva1 A 
.print op v(1) i(I1)
.op

.end
