* test for substitution
.options dollar_as_spice_comment

v1 n1 0 dc 1
.get     $PWD/ginclude/lib_file4.ckt
v2 n2 0 dc 2
.list
#.print op v(n*)
#.op
.end
